// Async fifo DUT
