// fifomem
