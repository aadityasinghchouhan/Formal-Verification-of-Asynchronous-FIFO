// rptr_empty
